module main (output  LED1, output  LED0);
assign LED1 = 1'b1;
assign LED0 = 1'b1;
endmodule

