module main (output  LED0, output  LED1);
assign LED0 = 1'b1;
assign LED1 = 1'b1;
endmodule

