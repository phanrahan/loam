module main (output  D1);
assign D1 = 1'b1;
endmodule

