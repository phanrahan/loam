module Register4 (input [3:0] I, output [3:0] O, input  CLK);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
SB_DFF inst0 (.C(CLK), .D(I[0]), .Q(inst0_Q));
SB_DFF inst1 (.C(CLK), .D(I[1]), .Q(inst1_Q));
SB_DFF inst2 (.C(CLK), .D(I[2]), .Q(inst2_Q));
SB_DFF inst3 (.C(CLK), .D(I[3]), .Q(inst3_Q));
assign O = {inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module main (input [4:0] J1, output [3:0] J3, input  CLKIN);
wire [3:0] inst0_O;
wire  inst1_out;
Register4 inst0 (.O(inst0_O), .CLK(inst1_out));
coreir_bitand inst1 (.in0(CLKIN), .in1(J1[4]), .out(inst1_out));
assign J3 = inst0_O;
endmodule

