module main (input [7:0] J1, output [7:0] J3);
assign J3 = J1;
endmodule

