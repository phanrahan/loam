module main (output [1:0] LED);
assign LED = {1'b0,1'b1};
endmodule

