module main (input  J1, output  J3);
assign J3 = J1;
endmodule

