module main (input  PIN4, output  PIN5);
assign PIN5 = PIN4;
endmodule

