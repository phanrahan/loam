module main (output  LED0, output  LED1, input  SWITCH0, input  SWITCH1);
assign LED0 = SWITCH0;
assign LED1 = SWITCH1;
endmodule

