module main (output  D5);
assign D5 = 1'b1;
endmodule

