module main (output [6:0] Digit0, output [6:0] Digit1);
assign Digit0 = {1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
assign Digit1 = {1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
endmodule

