module XOr3 (input [2:0] I, output  O);
wire  inst0_O;
LUT3 #(.INIT(8'h96)) inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .O(inst0_O));
assign O = inst0_O;
endmodule

module And2 (input [1:0] I, output  O);
wire  inst0_O;
LUT2 #(.INIT(4'h8)) inst0 (.I0(I[0]), .I1(I[1]), .O(inst0_O));
assign O = inst0_O;
endmodule

module Or3 (input [2:0] I, output  O);
wire  inst0_O;
LUT3 #(.INIT(8'h01)) inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .O(inst0_O));
assign O = inst0_O;
endmodule

module Op (input  I0, input  I1, input  I2, output  O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
And2 inst0 (.I({I1,I0}), .O(inst0_O));
And2 inst1 (.I({I2,I1}), .O(inst1_O));
And2 inst2 (.I({I0,I2}), .O(inst2_O));
Or3 inst3 (.I({inst2_O,inst1_O,inst0_O}), .O(inst3_O));
assign O = inst3_O;
endmodule

module PopCount128 (input [127:0] I, output [7:0] O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
wire  inst8_O;
wire  inst9_O;
wire  inst10_O;
wire  inst11_O;
wire  inst12_O;
wire  inst13_O;
wire  inst14_O;
wire  inst15_O;
wire  inst16_O;
wire  inst17_O;
wire  inst18_O;
wire  inst19_O;
wire  inst20_O;
wire  inst21_O;
wire  inst22_O;
wire  inst23_O;
wire  inst24_O;
wire  inst25_O;
wire  inst26_O;
wire  inst27_O;
wire  inst28_O;
wire  inst29_O;
wire  inst30_O;
wire  inst31_O;
wire  inst32_O;
wire  inst33_O;
wire  inst34_O;
wire  inst35_O;
wire  inst36_O;
wire  inst37_O;
wire  inst38_O;
wire  inst39_O;
wire  inst40_O;
wire  inst41_O;
wire  inst42_O;
wire  inst43_O;
wire  inst44_O;
wire  inst45_O;
wire  inst46_O;
wire  inst47_O;
wire  inst48_O;
wire  inst49_O;
wire  inst50_O;
wire  inst51_O;
wire  inst52_O;
wire  inst53_O;
wire  inst54_O;
wire  inst55_O;
wire  inst56_O;
wire  inst57_O;
wire  inst58_O;
wire  inst59_O;
wire  inst60_O;
wire  inst61_O;
wire  inst62_O;
wire  inst63_O;
wire  inst64_O;
wire  inst65_O;
wire  inst66_O;
wire  inst67_O;
wire  inst68_O;
wire  inst69_O;
wire  inst70_O;
wire  inst71_O;
wire  inst72_O;
wire  inst73_O;
wire  inst74_O;
wire  inst75_O;
wire  inst76_O;
wire  inst77_O;
wire  inst78_O;
wire  inst79_O;
wire  inst80_O;
wire  inst81_O;
wire  inst82_O;
wire  inst83_O;
wire  inst84_O;
wire  inst85_O;
wire  inst86_O;
wire  inst87_O;
wire  inst88_O;
wire  inst89_O;
wire  inst90_O;
wire  inst91_O;
wire  inst92_O;
wire  inst93_O;
wire  inst94_O;
wire  inst95_O;
wire  inst96_O;
wire  inst97_O;
wire  inst98_O;
wire  inst99_O;
wire  inst100_O;
wire  inst101_O;
wire  inst102_O;
wire  inst103_O;
wire  inst104_O;
wire  inst105_O;
wire  inst106_O;
wire  inst107_O;
wire  inst108_O;
wire  inst109_O;
wire  inst110_O;
wire  inst111_O;
wire  inst112_O;
wire  inst113_O;
wire  inst114_O;
wire  inst115_O;
wire  inst116_O;
wire  inst117_O;
wire  inst118_O;
wire  inst119_O;
wire  inst120_O;
wire  inst121_O;
wire  inst122_O;
wire  inst123_O;
wire  inst124_O;
wire  inst125_O;
wire  inst126_O;
wire  inst127_O;
wire  inst128_O;
wire  inst129_O;
wire  inst130_O;
wire  inst131_O;
wire  inst132_O;
wire  inst133_O;
wire  inst134_O;
wire  inst135_O;
wire  inst136_O;
wire  inst137_O;
wire  inst138_O;
wire  inst139_O;
wire  inst140_O;
wire  inst141_O;
wire  inst142_O;
wire  inst143_O;
wire  inst144_O;
wire  inst145_O;
wire  inst146_O;
wire  inst147_O;
wire  inst148_O;
wire  inst149_O;
wire  inst150_O;
wire  inst151_O;
wire  inst152_O;
wire  inst153_O;
wire  inst154_O;
wire  inst155_O;
wire  inst156_O;
wire  inst157_O;
wire  inst158_O;
wire  inst159_O;
wire  inst160_O;
wire  inst161_O;
wire  inst162_O;
wire  inst163_O;
wire  inst164_O;
wire  inst165_O;
wire  inst166_O;
wire  inst167_O;
wire  inst168_O;
wire  inst169_O;
wire  inst170_O;
wire  inst171_O;
wire  inst172_O;
wire  inst173_O;
wire  inst174_O;
wire  inst175_O;
wire  inst176_O;
wire  inst177_O;
wire  inst178_O;
wire  inst179_O;
wire  inst180_O;
wire  inst181_O;
wire  inst182_O;
wire  inst183_O;
wire  inst184_O;
wire  inst185_O;
wire  inst186_O;
wire  inst187_O;
wire  inst188_O;
wire  inst189_O;
wire  inst190_O;
wire  inst191_O;
wire  inst192_O;
wire  inst193_O;
wire  inst194_O;
wire  inst195_O;
wire  inst196_O;
wire  inst197_O;
wire  inst198_O;
wire  inst199_O;
wire  inst200_O;
wire  inst201_O;
wire  inst202_O;
wire  inst203_O;
wire  inst204_O;
wire  inst205_O;
wire  inst206_O;
wire  inst207_O;
wire  inst208_O;
wire  inst209_O;
wire  inst210_O;
wire  inst211_O;
wire  inst212_O;
wire  inst213_O;
wire  inst214_O;
wire  inst215_O;
wire  inst216_O;
wire  inst217_O;
wire  inst218_O;
wire  inst219_O;
wire  inst220_O;
wire  inst221_O;
wire  inst222_O;
wire  inst223_O;
wire  inst224_O;
wire  inst225_O;
wire  inst226_O;
wire  inst227_O;
wire  inst228_O;
wire  inst229_O;
wire  inst230_O;
wire  inst231_O;
wire  inst232_O;
wire  inst233_O;
wire  inst234_O;
wire  inst235_O;
wire  inst236_O;
wire  inst237_O;
wire  inst238_O;
wire  inst239_O;
wire  inst240_O;
wire  inst241_O;
wire  inst242_O;
wire  inst243_O;
wire  inst244_O;
wire  inst245_O;
wire  inst246_O;
wire  inst247_O;
wire  inst248_O;
wire  inst249_O;
wire  inst250_O;
wire  inst251_O;
wire  inst252_O;
wire  inst253_O;
XOr3 inst0 (.I({I[2],I[1],I[0]}), .O(inst0_O));
Op inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .O(inst1_O));
XOr3 inst2 (.I({I[5],I[4],I[3]}), .O(inst2_O));
Op inst3 (.I0(I[3]), .I1(I[4]), .I2(I[5]), .O(inst3_O));
XOr3 inst4 (.I({I[8],I[7],I[6]}), .O(inst4_O));
Op inst5 (.I0(I[6]), .I1(I[7]), .I2(I[8]), .O(inst5_O));
XOr3 inst6 (.I({I[11],I[10],I[9]}), .O(inst6_O));
Op inst7 (.I0(I[9]), .I1(I[10]), .I2(I[11]), .O(inst7_O));
XOr3 inst8 (.I({I[14],I[13],I[12]}), .O(inst8_O));
Op inst9 (.I0(I[12]), .I1(I[13]), .I2(I[14]), .O(inst9_O));
XOr3 inst10 (.I({I[17],I[16],I[15]}), .O(inst10_O));
Op inst11 (.I0(I[15]), .I1(I[16]), .I2(I[17]), .O(inst11_O));
XOr3 inst12 (.I({I[20],I[19],I[18]}), .O(inst12_O));
Op inst13 (.I0(I[18]), .I1(I[19]), .I2(I[20]), .O(inst13_O));
XOr3 inst14 (.I({I[23],I[22],I[21]}), .O(inst14_O));
Op inst15 (.I0(I[21]), .I1(I[22]), .I2(I[23]), .O(inst15_O));
XOr3 inst16 (.I({I[26],I[25],I[24]}), .O(inst16_O));
Op inst17 (.I0(I[24]), .I1(I[25]), .I2(I[26]), .O(inst17_O));
XOr3 inst18 (.I({I[29],I[28],I[27]}), .O(inst18_O));
Op inst19 (.I0(I[27]), .I1(I[28]), .I2(I[29]), .O(inst19_O));
XOr3 inst20 (.I({I[32],I[31],I[30]}), .O(inst20_O));
Op inst21 (.I0(I[30]), .I1(I[31]), .I2(I[32]), .O(inst21_O));
XOr3 inst22 (.I({I[35],I[34],I[33]}), .O(inst22_O));
Op inst23 (.I0(I[33]), .I1(I[34]), .I2(I[35]), .O(inst23_O));
XOr3 inst24 (.I({I[38],I[37],I[36]}), .O(inst24_O));
Op inst25 (.I0(I[36]), .I1(I[37]), .I2(I[38]), .O(inst25_O));
XOr3 inst26 (.I({I[41],I[40],I[39]}), .O(inst26_O));
Op inst27 (.I0(I[39]), .I1(I[40]), .I2(I[41]), .O(inst27_O));
XOr3 inst28 (.I({I[44],I[43],I[42]}), .O(inst28_O));
Op inst29 (.I0(I[42]), .I1(I[43]), .I2(I[44]), .O(inst29_O));
XOr3 inst30 (.I({I[47],I[46],I[45]}), .O(inst30_O));
Op inst31 (.I0(I[45]), .I1(I[46]), .I2(I[47]), .O(inst31_O));
XOr3 inst32 (.I({I[50],I[49],I[48]}), .O(inst32_O));
Op inst33 (.I0(I[48]), .I1(I[49]), .I2(I[50]), .O(inst33_O));
XOr3 inst34 (.I({I[53],I[52],I[51]}), .O(inst34_O));
Op inst35 (.I0(I[51]), .I1(I[52]), .I2(I[53]), .O(inst35_O));
XOr3 inst36 (.I({I[56],I[55],I[54]}), .O(inst36_O));
Op inst37 (.I0(I[54]), .I1(I[55]), .I2(I[56]), .O(inst37_O));
XOr3 inst38 (.I({I[59],I[58],I[57]}), .O(inst38_O));
Op inst39 (.I0(I[57]), .I1(I[58]), .I2(I[59]), .O(inst39_O));
XOr3 inst40 (.I({I[62],I[61],I[60]}), .O(inst40_O));
Op inst41 (.I0(I[60]), .I1(I[61]), .I2(I[62]), .O(inst41_O));
XOr3 inst42 (.I({I[65],I[64],I[63]}), .O(inst42_O));
Op inst43 (.I0(I[63]), .I1(I[64]), .I2(I[65]), .O(inst43_O));
XOr3 inst44 (.I({I[68],I[67],I[66]}), .O(inst44_O));
Op inst45 (.I0(I[66]), .I1(I[67]), .I2(I[68]), .O(inst45_O));
XOr3 inst46 (.I({I[71],I[70],I[69]}), .O(inst46_O));
Op inst47 (.I0(I[69]), .I1(I[70]), .I2(I[71]), .O(inst47_O));
XOr3 inst48 (.I({I[74],I[73],I[72]}), .O(inst48_O));
Op inst49 (.I0(I[72]), .I1(I[73]), .I2(I[74]), .O(inst49_O));
XOr3 inst50 (.I({I[77],I[76],I[75]}), .O(inst50_O));
Op inst51 (.I0(I[75]), .I1(I[76]), .I2(I[77]), .O(inst51_O));
XOr3 inst52 (.I({I[80],I[79],I[78]}), .O(inst52_O));
Op inst53 (.I0(I[78]), .I1(I[79]), .I2(I[80]), .O(inst53_O));
XOr3 inst54 (.I({I[83],I[82],I[81]}), .O(inst54_O));
Op inst55 (.I0(I[81]), .I1(I[82]), .I2(I[83]), .O(inst55_O));
XOr3 inst56 (.I({I[86],I[85],I[84]}), .O(inst56_O));
Op inst57 (.I0(I[84]), .I1(I[85]), .I2(I[86]), .O(inst57_O));
XOr3 inst58 (.I({I[89],I[88],I[87]}), .O(inst58_O));
Op inst59 (.I0(I[87]), .I1(I[88]), .I2(I[89]), .O(inst59_O));
XOr3 inst60 (.I({I[92],I[91],I[90]}), .O(inst60_O));
Op inst61 (.I0(I[90]), .I1(I[91]), .I2(I[92]), .O(inst61_O));
XOr3 inst62 (.I({I[95],I[94],I[93]}), .O(inst62_O));
Op inst63 (.I0(I[93]), .I1(I[94]), .I2(I[95]), .O(inst63_O));
XOr3 inst64 (.I({I[98],I[97],I[96]}), .O(inst64_O));
Op inst65 (.I0(I[96]), .I1(I[97]), .I2(I[98]), .O(inst65_O));
XOr3 inst66 (.I({I[101],I[100],I[99]}), .O(inst66_O));
Op inst67 (.I0(I[99]), .I1(I[100]), .I2(I[101]), .O(inst67_O));
XOr3 inst68 (.I({I[104],I[103],I[102]}), .O(inst68_O));
Op inst69 (.I0(I[102]), .I1(I[103]), .I2(I[104]), .O(inst69_O));
XOr3 inst70 (.I({I[107],I[106],I[105]}), .O(inst70_O));
Op inst71 (.I0(I[105]), .I1(I[106]), .I2(I[107]), .O(inst71_O));
XOr3 inst72 (.I({I[110],I[109],I[108]}), .O(inst72_O));
Op inst73 (.I0(I[108]), .I1(I[109]), .I2(I[110]), .O(inst73_O));
XOr3 inst74 (.I({I[113],I[112],I[111]}), .O(inst74_O));
Op inst75 (.I0(I[111]), .I1(I[112]), .I2(I[113]), .O(inst75_O));
XOr3 inst76 (.I({I[116],I[115],I[114]}), .O(inst76_O));
Op inst77 (.I0(I[114]), .I1(I[115]), .I2(I[116]), .O(inst77_O));
XOr3 inst78 (.I({I[119],I[118],I[117]}), .O(inst78_O));
Op inst79 (.I0(I[117]), .I1(I[118]), .I2(I[119]), .O(inst79_O));
XOr3 inst80 (.I({I[122],I[121],I[120]}), .O(inst80_O));
Op inst81 (.I0(I[120]), .I1(I[121]), .I2(I[122]), .O(inst81_O));
XOr3 inst82 (.I({I[125],I[124],I[123]}), .O(inst82_O));
Op inst83 (.I0(I[123]), .I1(I[124]), .I2(I[125]), .O(inst83_O));
XOr3 inst84 (.I({inst4_O,inst2_O,inst0_O}), .O(inst84_O));
Op inst85 (.I0(inst0_O), .I1(inst2_O), .I2(inst4_O), .O(inst85_O));
XOr3 inst86 (.I({inst10_O,inst8_O,inst6_O}), .O(inst86_O));
Op inst87 (.I0(inst6_O), .I1(inst8_O), .I2(inst10_O), .O(inst87_O));
XOr3 inst88 (.I({inst16_O,inst14_O,inst12_O}), .O(inst88_O));
Op inst89 (.I0(inst12_O), .I1(inst14_O), .I2(inst16_O), .O(inst89_O));
XOr3 inst90 (.I({inst22_O,inst20_O,inst18_O}), .O(inst90_O));
Op inst91 (.I0(inst18_O), .I1(inst20_O), .I2(inst22_O), .O(inst91_O));
XOr3 inst92 (.I({inst28_O,inst26_O,inst24_O}), .O(inst92_O));
Op inst93 (.I0(inst24_O), .I1(inst26_O), .I2(inst28_O), .O(inst93_O));
XOr3 inst94 (.I({inst34_O,inst32_O,inst30_O}), .O(inst94_O));
Op inst95 (.I0(inst30_O), .I1(inst32_O), .I2(inst34_O), .O(inst95_O));
XOr3 inst96 (.I({inst40_O,inst38_O,inst36_O}), .O(inst96_O));
Op inst97 (.I0(inst36_O), .I1(inst38_O), .I2(inst40_O), .O(inst97_O));
XOr3 inst98 (.I({inst46_O,inst44_O,inst42_O}), .O(inst98_O));
Op inst99 (.I0(inst42_O), .I1(inst44_O), .I2(inst46_O), .O(inst99_O));
XOr3 inst100 (.I({inst52_O,inst50_O,inst48_O}), .O(inst100_O));
Op inst101 (.I0(inst48_O), .I1(inst50_O), .I2(inst52_O), .O(inst101_O));
XOr3 inst102 (.I({inst58_O,inst56_O,inst54_O}), .O(inst102_O));
Op inst103 (.I0(inst54_O), .I1(inst56_O), .I2(inst58_O), .O(inst103_O));
XOr3 inst104 (.I({inst64_O,inst62_O,inst60_O}), .O(inst104_O));
Op inst105 (.I0(inst60_O), .I1(inst62_O), .I2(inst64_O), .O(inst105_O));
XOr3 inst106 (.I({inst70_O,inst68_O,inst66_O}), .O(inst106_O));
Op inst107 (.I0(inst66_O), .I1(inst68_O), .I2(inst70_O), .O(inst107_O));
XOr3 inst108 (.I({inst76_O,inst74_O,inst72_O}), .O(inst108_O));
Op inst109 (.I0(inst72_O), .I1(inst74_O), .I2(inst76_O), .O(inst109_O));
XOr3 inst110 (.I({inst82_O,inst80_O,inst78_O}), .O(inst110_O));
Op inst111 (.I0(inst78_O), .I1(inst80_O), .I2(inst82_O), .O(inst111_O));
XOr3 inst112 (.I({inst5_O,inst3_O,inst1_O}), .O(inst112_O));
Op inst113 (.I0(inst1_O), .I1(inst3_O), .I2(inst5_O), .O(inst113_O));
XOr3 inst114 (.I({inst11_O,inst9_O,inst7_O}), .O(inst114_O));
Op inst115 (.I0(inst7_O), .I1(inst9_O), .I2(inst11_O), .O(inst115_O));
XOr3 inst116 (.I({inst17_O,inst15_O,inst13_O}), .O(inst116_O));
Op inst117 (.I0(inst13_O), .I1(inst15_O), .I2(inst17_O), .O(inst117_O));
XOr3 inst118 (.I({inst23_O,inst21_O,inst19_O}), .O(inst118_O));
Op inst119 (.I0(inst19_O), .I1(inst21_O), .I2(inst23_O), .O(inst119_O));
XOr3 inst120 (.I({inst29_O,inst27_O,inst25_O}), .O(inst120_O));
Op inst121 (.I0(inst25_O), .I1(inst27_O), .I2(inst29_O), .O(inst121_O));
XOr3 inst122 (.I({inst35_O,inst33_O,inst31_O}), .O(inst122_O));
Op inst123 (.I0(inst31_O), .I1(inst33_O), .I2(inst35_O), .O(inst123_O));
XOr3 inst124 (.I({inst41_O,inst39_O,inst37_O}), .O(inst124_O));
Op inst125 (.I0(inst37_O), .I1(inst39_O), .I2(inst41_O), .O(inst125_O));
XOr3 inst126 (.I({inst47_O,inst45_O,inst43_O}), .O(inst126_O));
Op inst127 (.I0(inst43_O), .I1(inst45_O), .I2(inst47_O), .O(inst127_O));
XOr3 inst128 (.I({inst53_O,inst51_O,inst49_O}), .O(inst128_O));
Op inst129 (.I0(inst49_O), .I1(inst51_O), .I2(inst53_O), .O(inst129_O));
XOr3 inst130 (.I({inst59_O,inst57_O,inst55_O}), .O(inst130_O));
Op inst131 (.I0(inst55_O), .I1(inst57_O), .I2(inst59_O), .O(inst131_O));
XOr3 inst132 (.I({inst65_O,inst63_O,inst61_O}), .O(inst132_O));
Op inst133 (.I0(inst61_O), .I1(inst63_O), .I2(inst65_O), .O(inst133_O));
XOr3 inst134 (.I({inst71_O,inst69_O,inst67_O}), .O(inst134_O));
Op inst135 (.I0(inst67_O), .I1(inst69_O), .I2(inst71_O), .O(inst135_O));
XOr3 inst136 (.I({inst77_O,inst75_O,inst73_O}), .O(inst136_O));
Op inst137 (.I0(inst73_O), .I1(inst75_O), .I2(inst77_O), .O(inst137_O));
XOr3 inst138 (.I({inst83_O,inst81_O,inst79_O}), .O(inst138_O));
Op inst139 (.I0(inst79_O), .I1(inst81_O), .I2(inst83_O), .O(inst139_O));
XOr3 inst140 (.I({inst88_O,inst86_O,inst84_O}), .O(inst140_O));
Op inst141 (.I0(inst84_O), .I1(inst86_O), .I2(inst88_O), .O(inst141_O));
XOr3 inst142 (.I({inst94_O,inst92_O,inst90_O}), .O(inst142_O));
Op inst143 (.I0(inst90_O), .I1(inst92_O), .I2(inst94_O), .O(inst143_O));
XOr3 inst144 (.I({inst100_O,inst98_O,inst96_O}), .O(inst144_O));
Op inst145 (.I0(inst96_O), .I1(inst98_O), .I2(inst100_O), .O(inst145_O));
XOr3 inst146 (.I({inst106_O,inst104_O,inst102_O}), .O(inst146_O));
Op inst147 (.I0(inst102_O), .I1(inst104_O), .I2(inst106_O), .O(inst147_O));
XOr3 inst148 (.I({I[126],inst110_O,inst108_O}), .O(inst148_O));
Op inst149 (.I0(inst108_O), .I1(inst110_O), .I2(I[126]), .O(inst149_O));
XOr3 inst150 (.I({inst116_O,inst114_O,inst112_O}), .O(inst150_O));
Op inst151 (.I0(inst112_O), .I1(inst114_O), .I2(inst116_O), .O(inst151_O));
XOr3 inst152 (.I({inst122_O,inst120_O,inst118_O}), .O(inst152_O));
Op inst153 (.I0(inst118_O), .I1(inst120_O), .I2(inst122_O), .O(inst153_O));
XOr3 inst154 (.I({inst128_O,inst126_O,inst124_O}), .O(inst154_O));
Op inst155 (.I0(inst124_O), .I1(inst126_O), .I2(inst128_O), .O(inst155_O));
XOr3 inst156 (.I({inst134_O,inst132_O,inst130_O}), .O(inst156_O));
Op inst157 (.I0(inst130_O), .I1(inst132_O), .I2(inst134_O), .O(inst157_O));
XOr3 inst158 (.I({inst85_O,inst138_O,inst136_O}), .O(inst158_O));
Op inst159 (.I0(inst136_O), .I1(inst138_O), .I2(inst85_O), .O(inst159_O));
XOr3 inst160 (.I({inst91_O,inst89_O,inst87_O}), .O(inst160_O));
Op inst161 (.I0(inst87_O), .I1(inst89_O), .I2(inst91_O), .O(inst161_O));
XOr3 inst162 (.I({inst97_O,inst95_O,inst93_O}), .O(inst162_O));
Op inst163 (.I0(inst93_O), .I1(inst95_O), .I2(inst97_O), .O(inst163_O));
XOr3 inst164 (.I({inst103_O,inst101_O,inst99_O}), .O(inst164_O));
Op inst165 (.I0(inst99_O), .I1(inst101_O), .I2(inst103_O), .O(inst165_O));
XOr3 inst166 (.I({inst109_O,inst107_O,inst105_O}), .O(inst166_O));
Op inst167 (.I0(inst105_O), .I1(inst107_O), .I2(inst109_O), .O(inst167_O));
XOr3 inst168 (.I({inst117_O,inst115_O,inst113_O}), .O(inst168_O));
Op inst169 (.I0(inst113_O), .I1(inst115_O), .I2(inst117_O), .O(inst169_O));
XOr3 inst170 (.I({inst123_O,inst121_O,inst119_O}), .O(inst170_O));
Op inst171 (.I0(inst119_O), .I1(inst121_O), .I2(inst123_O), .O(inst171_O));
XOr3 inst172 (.I({inst129_O,inst127_O,inst125_O}), .O(inst172_O));
Op inst173 (.I0(inst125_O), .I1(inst127_O), .I2(inst129_O), .O(inst173_O));
XOr3 inst174 (.I({inst135_O,inst133_O,inst131_O}), .O(inst174_O));
Op inst175 (.I0(inst131_O), .I1(inst133_O), .I2(inst135_O), .O(inst175_O));
XOr3 inst176 (.I({inst144_O,inst142_O,inst140_O}), .O(inst176_O));
Op inst177 (.I0(inst140_O), .I1(inst142_O), .I2(inst144_O), .O(inst177_O));
XOr3 inst178 (.I({I[127],inst148_O,inst146_O}), .O(inst178_O));
Op inst179 (.I0(inst146_O), .I1(inst148_O), .I2(I[127]), .O(inst179_O));
XOr3 inst180 (.I({inst154_O,inst152_O,inst150_O}), .O(inst180_O));
Op inst181 (.I0(inst150_O), .I1(inst152_O), .I2(inst154_O), .O(inst181_O));
XOr3 inst182 (.I({inst160_O,inst158_O,inst156_O}), .O(inst182_O));
Op inst183 (.I0(inst156_O), .I1(inst158_O), .I2(inst160_O), .O(inst183_O));
XOr3 inst184 (.I({inst166_O,inst164_O,inst162_O}), .O(inst184_O));
Op inst185 (.I0(inst162_O), .I1(inst164_O), .I2(inst166_O), .O(inst185_O));
XOr3 inst186 (.I({inst143_O,inst141_O,inst111_O}), .O(inst186_O));
Op inst187 (.I0(inst111_O), .I1(inst141_O), .I2(inst143_O), .O(inst187_O));
XOr3 inst188 (.I({inst149_O,inst147_O,inst145_O}), .O(inst188_O));
Op inst189 (.I0(inst145_O), .I1(inst147_O), .I2(inst149_O), .O(inst189_O));
XOr3 inst190 (.I({inst172_O,inst170_O,inst168_O}), .O(inst190_O));
Op inst191 (.I0(inst168_O), .I1(inst170_O), .I2(inst172_O), .O(inst191_O));
XOr3 inst192 (.I({inst139_O,inst137_O,inst174_O}), .O(inst192_O));
Op inst193 (.I0(inst174_O), .I1(inst137_O), .I2(inst139_O), .O(inst193_O));
XOr3 inst194 (.I({inst155_O,inst153_O,inst151_O}), .O(inst194_O));
Op inst195 (.I0(inst151_O), .I1(inst153_O), .I2(inst155_O), .O(inst195_O));
XOr3 inst196 (.I({inst161_O,inst159_O,inst157_O}), .O(inst196_O));
Op inst197 (.I0(inst157_O), .I1(inst159_O), .I2(inst161_O), .O(inst197_O));
XOr3 inst198 (.I({inst167_O,inst165_O,inst163_O}), .O(inst198_O));
Op inst199 (.I0(inst163_O), .I1(inst165_O), .I2(inst167_O), .O(inst199_O));
XOr3 inst200 (.I({inst173_O,inst171_O,inst169_O}), .O(inst200_O));
Op inst201 (.I0(inst169_O), .I1(inst171_O), .I2(inst173_O), .O(inst201_O));
XOr3 inst202 (.I({inst184_O,inst182_O,inst180_O}), .O(inst202_O));
Op inst203 (.I0(inst180_O), .I1(inst182_O), .I2(inst184_O), .O(inst203_O));
XOr3 inst204 (.I({inst177_O,inst188_O,inst186_O}), .O(inst204_O));
Op inst205 (.I0(inst186_O), .I1(inst188_O), .I2(inst177_O), .O(inst205_O));
XOr3 inst206 (.I({inst194_O,inst192_O,inst190_O}), .O(inst206_O));
Op inst207 (.I0(inst190_O), .I1(inst192_O), .I2(inst194_O), .O(inst207_O));
XOr3 inst208 (.I({inst181_O,inst198_O,inst196_O}), .O(inst208_O));
Op inst209 (.I0(inst196_O), .I1(inst198_O), .I2(inst181_O), .O(inst209_O));
XOr3 inst210 (.I({inst187_O,inst185_O,inst183_O}), .O(inst210_O));
Op inst211 (.I0(inst183_O), .I1(inst185_O), .I2(inst187_O), .O(inst211_O));
XOr3 inst212 (.I({inst191_O,inst175_O,inst200_O}), .O(inst212_O));
Op inst213 (.I0(inst200_O), .I1(inst175_O), .I2(inst191_O), .O(inst213_O));
XOr3 inst214 (.I({inst197_O,inst195_O,inst193_O}), .O(inst214_O));
Op inst215 (.I0(inst193_O), .I1(inst195_O), .I2(inst197_O), .O(inst215_O));
XOr3 inst216 (.I({inst179_O,inst204_O,inst202_O}), .O(inst216_O));
Op inst217 (.I0(inst202_O), .I1(inst204_O), .I2(inst179_O), .O(inst217_O));
XOr3 inst218 (.I({inst210_O,inst208_O,inst206_O}), .O(inst218_O));
Op inst219 (.I0(inst206_O), .I1(inst208_O), .I2(inst210_O), .O(inst219_O));
XOr3 inst220 (.I({inst205_O,inst203_O,inst189_O}), .O(inst220_O));
Op inst221 (.I0(inst189_O), .I1(inst203_O), .I2(inst205_O), .O(inst221_O));
XOr3 inst222 (.I({inst199_O,inst214_O,inst212_O}), .O(inst222_O));
Op inst223 (.I0(inst212_O), .I1(inst214_O), .I2(inst199_O), .O(inst223_O));
XOr3 inst224 (.I({inst211_O,inst209_O,inst207_O}), .O(inst224_O));
Op inst225 (.I0(inst207_O), .I1(inst209_O), .I2(inst211_O), .O(inst225_O));
XOr3 inst226 (.I({inst215_O,inst213_O,inst201_O}), .O(inst226_O));
Op inst227 (.I0(inst201_O), .I1(inst213_O), .I2(inst215_O), .O(inst227_O));
XOr3 inst228 (.I({inst217_O,inst220_O,inst218_O}), .O(inst228_O));
Op inst229 (.I0(inst218_O), .I1(inst220_O), .I2(inst217_O), .O(inst229_O));
XOr3 inst230 (.I({inst219_O,inst224_O,inst222_O}), .O(inst230_O));
Op inst231 (.I0(inst222_O), .I1(inst224_O), .I2(inst219_O), .O(inst231_O));
XOr3 inst232 (.I({inst225_O,inst223_O,inst226_O}), .O(inst232_O));
Op inst233 (.I0(inst226_O), .I1(inst223_O), .I2(inst225_O), .O(inst233_O));
XOr3 inst234 (.I({inst229_O,inst221_O,inst230_O}), .O(inst234_O));
Op inst235 (.I0(inst230_O), .I1(inst221_O), .I2(inst229_O), .O(inst235_O));
XOr3 inst236 (.I({inst235_O,inst231_O,inst232_O}), .O(inst236_O));
Op inst237 (.I0(inst232_O), .I1(inst231_O), .I2(inst235_O), .O(inst237_O));
XOr3 inst238 (.I({inst237_O,inst233_O,inst227_O}), .O(inst238_O));
Op inst239 (.I0(inst227_O), .I1(inst233_O), .I2(inst237_O), .O(inst239_O));
XOr3 inst240 (.I({1'b0,inst178_O,inst176_O}), .O(inst240_O));
Op inst241 (.I0(inst176_O), .I1(inst178_O), .I2(1'b0), .O(inst241_O));
XOr3 inst242 (.I({1'b0,inst241_O,inst216_O}), .O(inst242_O));
Op inst243 (.I0(inst216_O), .I1(inst241_O), .I2(1'b0), .O(inst243_O));
XOr3 inst244 (.I({1'b0,inst243_O,inst228_O}), .O(inst244_O));
Op inst245 (.I0(inst228_O), .I1(inst243_O), .I2(1'b0), .O(inst245_O));
XOr3 inst246 (.I({1'b0,inst245_O,inst234_O}), .O(inst246_O));
Op inst247 (.I0(inst234_O), .I1(inst245_O), .I2(1'b0), .O(inst247_O));
XOr3 inst248 (.I({1'b0,inst247_O,inst236_O}), .O(inst248_O));
Op inst249 (.I0(inst236_O), .I1(inst247_O), .I2(1'b0), .O(inst249_O));
XOr3 inst250 (.I({1'b0,inst249_O,inst238_O}), .O(inst250_O));
Op inst251 (.I0(inst238_O), .I1(inst249_O), .I2(1'b0), .O(inst251_O));
XOr3 inst252 (.I({1'b0,inst251_O,inst239_O}), .O(inst252_O));
Op inst253 (.I0(inst239_O), .I1(inst251_O), .I2(1'b0), .O(inst253_O));
assign O = {inst253_O,inst252_O,inst250_O,inst248_O,inst246_O,inst244_O,inst242_O,inst240_O};
endmodule

module main (input [7:0] SWITCH, output [7:0] LED);
wire [7:0] inst0_O;
PopCount128 inst0 (.I({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,SWITCH[7],SWITCH[6],SWITCH[5],SWITCH[4],SWITCH[3],SWITCH[2],SWITCH[1],SWITCH[0]}), .O(inst0_O));
assign LED = inst0_O;
endmodule

