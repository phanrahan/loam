module main (output [0:0] LED);
assign LED = {1'b1};
endmodule

