module main (output  LED_R);
assign LED_R = 1'b1;
endmodule

