module main (output  D1, output  D2);
assign D1 = 1'b1;
assign D2 = 1'b1;
endmodule

