module main (input  B1, output  D1);
assign D1 = B1;
endmodule

