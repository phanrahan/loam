module main (input [3:0] J1i, output [3:0] J1o, input  CLKIN);
assign J1o = J1i;
endmodule

