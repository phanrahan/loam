module Decode8 (input [7:0] I, output  O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
wire  inst8_O;
wire  inst9_O;
wire  inst10_O;
wire  inst11_O;
wire  inst12_O;
wire  inst13_O;
wire  inst14_O;
wire  inst15_O;
wire  inst16_O;
wire  inst17_O;
wire  inst18_O;
wire  inst19_O;
wire  inst20_O;
wire  inst21_O;
wire  inst22_O;
wire  inst23_O;
wire  inst24_O;
wire  inst25_O;
wire  inst26_O;
wire  inst27_O;
wire  inst28_O;
wire  inst29_O;
wire  inst30_O;
LUT4 #(.INIT(16'h0001)) inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst0_O));
LUT4 #(.INIT(16'h0000)) inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst1_O));
MUXF5 inst2 (.I0(inst0_O), .I1(inst1_O), .S(I[4]), .O(inst2_O));
LUT4 #(.INIT(16'h0000)) inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst3_O));
LUT4 #(.INIT(16'h0000)) inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst4_O));
MUXF5 inst5 (.I0(inst3_O), .I1(inst4_O), .S(I[4]), .O(inst5_O));
MUXF6 inst6 (.I0(inst2_O), .I1(inst5_O), .S(I[5]), .O(inst6_O));
LUT4 #(.INIT(16'h0000)) inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst7_O));
LUT4 #(.INIT(16'h0000)) inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst8_O));
MUXF5 inst9 (.I0(inst7_O), .I1(inst8_O), .S(I[4]), .O(inst9_O));
LUT4 #(.INIT(16'h0000)) inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst10_O));
LUT4 #(.INIT(16'h0000)) inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst11_O));
MUXF5 inst12 (.I0(inst10_O), .I1(inst11_O), .S(I[4]), .O(inst12_O));
MUXF6 inst13 (.I0(inst9_O), .I1(inst12_O), .S(I[5]), .O(inst13_O));
MUXF7 inst14 (.I0(inst6_O), .I1(inst13_O), .S(I[6]), .O(inst14_O));
LUT4 #(.INIT(16'h0000)) inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst15_O));
LUT4 #(.INIT(16'h0000)) inst16 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst16_O));
MUXF5 inst17 (.I0(inst15_O), .I1(inst16_O), .S(I[4]), .O(inst17_O));
LUT4 #(.INIT(16'h0000)) inst18 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst18_O));
LUT4 #(.INIT(16'h0000)) inst19 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst19_O));
MUXF5 inst20 (.I0(inst18_O), .I1(inst19_O), .S(I[4]), .O(inst20_O));
MUXF6 inst21 (.I0(inst17_O), .I1(inst20_O), .S(I[5]), .O(inst21_O));
LUT4 #(.INIT(16'h0000)) inst22 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst22_O));
LUT4 #(.INIT(16'h0000)) inst23 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst23_O));
MUXF5 inst24 (.I0(inst22_O), .I1(inst23_O), .S(I[4]), .O(inst24_O));
LUT4 #(.INIT(16'h0000)) inst25 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst25_O));
LUT4 #(.INIT(16'h0000)) inst26 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst26_O));
MUXF5 inst27 (.I0(inst25_O), .I1(inst26_O), .S(I[4]), .O(inst27_O));
MUXF6 inst28 (.I0(inst24_O), .I1(inst27_O), .S(I[5]), .O(inst28_O));
MUXF7 inst29 (.I0(inst21_O), .I1(inst28_O), .S(I[6]), .O(inst29_O));
MUXF8 inst30 (.I0(inst14_O), .I1(inst29_O), .S(I[7]), .O(inst30_O));
assign O = inst30_O;
endmodule

module main (input [7:0] SWITCH, output  LED);
wire  inst0_O;
Decode8 inst0 (.I(SWITCH), .O(inst0_O));
assign LED = inst0_O;
endmodule

