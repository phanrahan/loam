module main (output  LED1, output  LED0, input  SWITCH1, input  SWITCH0);
assign LED1 = SWITCH1;
assign LED0 = SWITCH0;
endmodule

