module main (output  PIN4);
assign PIN4 = 1'b1;
endmodule

