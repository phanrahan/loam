module main (output  PIN2, input  PIN3);
assign PIN2 = PIN3;
endmodule

