module Add32_cout (input [31:0] I0, input [31:0] I1, output [31:0] O, output  COUT);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
wire  inst8_O;
wire  inst9_O;
wire  inst10_O;
wire  inst11_O;
wire  inst12_O;
wire  inst13_O;
wire  inst14_O;
wire  inst15_O;
wire  inst16_O;
wire  inst17_O;
wire  inst18_O;
wire  inst19_O;
wire  inst20_O;
wire  inst21_O;
wire  inst22_O;
wire  inst23_O;
wire  inst24_O;
wire  inst25_O;
wire  inst26_O;
wire  inst27_O;
wire  inst28_O;
wire  inst29_O;
wire  inst30_O;
wire  inst31_O;
wire  inst32_O;
wire  inst33_O;
wire  inst34_O;
wire  inst35_O;
wire  inst36_O;
wire  inst37_O;
wire  inst38_O;
wire  inst39_O;
wire  inst40_O;
wire  inst41_O;
wire  inst42_O;
wire  inst43_O;
wire  inst44_O;
wire  inst45_O;
wire  inst46_O;
wire  inst47_O;
wire  inst48_O;
wire  inst49_O;
wire  inst50_O;
wire  inst51_O;
wire  inst52_O;
wire  inst53_O;
wire  inst54_O;
wire  inst55_O;
wire  inst56_O;
wire  inst57_O;
wire  inst58_O;
wire  inst59_O;
wire  inst60_O;
wire  inst61_O;
wire  inst62_O;
wire  inst63_O;
LUT2 #(.INIT(4'h6)) inst0 (.I0(I0[0]), .I1(I1[0]), .O(inst0_O));
MUXCY inst1 (.DI(I0[0]), .CI(1'b0), .S(inst0_O), .O(inst1_O));
LUT2 #(.INIT(4'h6)) inst2 (.I0(I0[1]), .I1(I1[1]), .O(inst2_O));
MUXCY inst3 (.DI(I0[1]), .CI(inst1_O), .S(inst2_O), .O(inst3_O));
LUT2 #(.INIT(4'h6)) inst4 (.I0(I0[2]), .I1(I1[2]), .O(inst4_O));
MUXCY inst5 (.DI(I0[2]), .CI(inst3_O), .S(inst4_O), .O(inst5_O));
LUT2 #(.INIT(4'h6)) inst6 (.I0(I0[3]), .I1(I1[3]), .O(inst6_O));
MUXCY inst7 (.DI(I0[3]), .CI(inst5_O), .S(inst6_O), .O(inst7_O));
LUT2 #(.INIT(4'h6)) inst8 (.I0(I0[4]), .I1(I1[4]), .O(inst8_O));
MUXCY inst9 (.DI(I0[4]), .CI(inst7_O), .S(inst8_O), .O(inst9_O));
LUT2 #(.INIT(4'h6)) inst10 (.I0(I0[5]), .I1(I1[5]), .O(inst10_O));
MUXCY inst11 (.DI(I0[5]), .CI(inst9_O), .S(inst10_O), .O(inst11_O));
LUT2 #(.INIT(4'h6)) inst12 (.I0(I0[6]), .I1(I1[6]), .O(inst12_O));
MUXCY inst13 (.DI(I0[6]), .CI(inst11_O), .S(inst12_O), .O(inst13_O));
LUT2 #(.INIT(4'h6)) inst14 (.I0(I0[7]), .I1(I1[7]), .O(inst14_O));
MUXCY inst15 (.DI(I0[7]), .CI(inst13_O), .S(inst14_O), .O(inst15_O));
LUT2 #(.INIT(4'h6)) inst16 (.I0(I0[8]), .I1(I1[8]), .O(inst16_O));
MUXCY inst17 (.DI(I0[8]), .CI(inst15_O), .S(inst16_O), .O(inst17_O));
LUT2 #(.INIT(4'h6)) inst18 (.I0(I0[9]), .I1(I1[9]), .O(inst18_O));
MUXCY inst19 (.DI(I0[9]), .CI(inst17_O), .S(inst18_O), .O(inst19_O));
LUT2 #(.INIT(4'h6)) inst20 (.I0(I0[10]), .I1(I1[10]), .O(inst20_O));
MUXCY inst21 (.DI(I0[10]), .CI(inst19_O), .S(inst20_O), .O(inst21_O));
LUT2 #(.INIT(4'h6)) inst22 (.I0(I0[11]), .I1(I1[11]), .O(inst22_O));
MUXCY inst23 (.DI(I0[11]), .CI(inst21_O), .S(inst22_O), .O(inst23_O));
LUT2 #(.INIT(4'h6)) inst24 (.I0(I0[12]), .I1(I1[12]), .O(inst24_O));
MUXCY inst25 (.DI(I0[12]), .CI(inst23_O), .S(inst24_O), .O(inst25_O));
LUT2 #(.INIT(4'h6)) inst26 (.I0(I0[13]), .I1(I1[13]), .O(inst26_O));
MUXCY inst27 (.DI(I0[13]), .CI(inst25_O), .S(inst26_O), .O(inst27_O));
LUT2 #(.INIT(4'h6)) inst28 (.I0(I0[14]), .I1(I1[14]), .O(inst28_O));
MUXCY inst29 (.DI(I0[14]), .CI(inst27_O), .S(inst28_O), .O(inst29_O));
LUT2 #(.INIT(4'h6)) inst30 (.I0(I0[15]), .I1(I1[15]), .O(inst30_O));
MUXCY inst31 (.DI(I0[15]), .CI(inst29_O), .S(inst30_O), .O(inst31_O));
LUT2 #(.INIT(4'h6)) inst32 (.I0(I0[16]), .I1(I1[16]), .O(inst32_O));
MUXCY inst33 (.DI(I0[16]), .CI(inst31_O), .S(inst32_O), .O(inst33_O));
LUT2 #(.INIT(4'h6)) inst34 (.I0(I0[17]), .I1(I1[17]), .O(inst34_O));
MUXCY inst35 (.DI(I0[17]), .CI(inst33_O), .S(inst34_O), .O(inst35_O));
LUT2 #(.INIT(4'h6)) inst36 (.I0(I0[18]), .I1(I1[18]), .O(inst36_O));
MUXCY inst37 (.DI(I0[18]), .CI(inst35_O), .S(inst36_O), .O(inst37_O));
LUT2 #(.INIT(4'h6)) inst38 (.I0(I0[19]), .I1(I1[19]), .O(inst38_O));
MUXCY inst39 (.DI(I0[19]), .CI(inst37_O), .S(inst38_O), .O(inst39_O));
LUT2 #(.INIT(4'h6)) inst40 (.I0(I0[20]), .I1(I1[20]), .O(inst40_O));
MUXCY inst41 (.DI(I0[20]), .CI(inst39_O), .S(inst40_O), .O(inst41_O));
LUT2 #(.INIT(4'h6)) inst42 (.I0(I0[21]), .I1(I1[21]), .O(inst42_O));
MUXCY inst43 (.DI(I0[21]), .CI(inst41_O), .S(inst42_O), .O(inst43_O));
LUT2 #(.INIT(4'h6)) inst44 (.I0(I0[22]), .I1(I1[22]), .O(inst44_O));
MUXCY inst45 (.DI(I0[22]), .CI(inst43_O), .S(inst44_O), .O(inst45_O));
LUT2 #(.INIT(4'h6)) inst46 (.I0(I0[23]), .I1(I1[23]), .O(inst46_O));
MUXCY inst47 (.DI(I0[23]), .CI(inst45_O), .S(inst46_O), .O(inst47_O));
LUT2 #(.INIT(4'h6)) inst48 (.I0(I0[24]), .I1(I1[24]), .O(inst48_O));
MUXCY inst49 (.DI(I0[24]), .CI(inst47_O), .S(inst48_O), .O(inst49_O));
LUT2 #(.INIT(4'h6)) inst50 (.I0(I0[25]), .I1(I1[25]), .O(inst50_O));
MUXCY inst51 (.DI(I0[25]), .CI(inst49_O), .S(inst50_O), .O(inst51_O));
LUT2 #(.INIT(4'h6)) inst52 (.I0(I0[26]), .I1(I1[26]), .O(inst52_O));
MUXCY inst53 (.DI(I0[26]), .CI(inst51_O), .S(inst52_O), .O(inst53_O));
LUT2 #(.INIT(4'h6)) inst54 (.I0(I0[27]), .I1(I1[27]), .O(inst54_O));
MUXCY inst55 (.DI(I0[27]), .CI(inst53_O), .S(inst54_O), .O(inst55_O));
LUT2 #(.INIT(4'h6)) inst56 (.I0(I0[28]), .I1(I1[28]), .O(inst56_O));
MUXCY inst57 (.DI(I0[28]), .CI(inst55_O), .S(inst56_O), .O(inst57_O));
LUT2 #(.INIT(4'h6)) inst58 (.I0(I0[29]), .I1(I1[29]), .O(inst58_O));
MUXCY inst59 (.DI(I0[29]), .CI(inst57_O), .S(inst58_O), .O(inst59_O));
LUT2 #(.INIT(4'h6)) inst60 (.I0(I0[30]), .I1(I1[30]), .O(inst60_O));
MUXCY inst61 (.DI(I0[30]), .CI(inst59_O), .S(inst60_O), .O(inst61_O));
LUT2 #(.INIT(4'h6)) inst62 (.I0(I0[31]), .I1(I1[31]), .O(inst62_O));
MUXCY inst63 (.DI(I0[31]), .CI(inst61_O), .S(inst62_O), .O(inst63_O));
assign O = {inst62_O,inst60_O,inst58_O,inst56_O,inst54_O,inst52_O,inst50_O,inst48_O,inst46_O,inst44_O,inst42_O,inst40_O,inst38_O,inst36_O,inst34_O,inst32_O,inst30_O,inst28_O,inst26_O,inst24_O,inst22_O,inst20_O,inst18_O,inst16_O,inst14_O,inst12_O,inst10_O,inst8_O,inst6_O,inst4_O,inst2_O,inst0_O};
assign COUT = inst63_O;
endmodule

module Register32 (input [31:0] I, output [31:0] O, input  CLK);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
wire  inst4_Q;
wire  inst5_Q;
wire  inst6_Q;
wire  inst7_Q;
wire  inst8_Q;
wire  inst9_Q;
wire  inst10_Q;
wire  inst11_Q;
wire  inst12_Q;
wire  inst13_Q;
wire  inst14_Q;
wire  inst15_Q;
wire  inst16_Q;
wire  inst17_Q;
wire  inst18_Q;
wire  inst19_Q;
wire  inst20_Q;
wire  inst21_Q;
wire  inst22_Q;
wire  inst23_Q;
wire  inst24_Q;
wire  inst25_Q;
wire  inst26_Q;
wire  inst27_Q;
wire  inst28_Q;
wire  inst29_Q;
wire  inst30_Q;
wire  inst31_Q;
FDRSE #(.INIT(1'h0)) inst0 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[0]), .Q(inst0_Q));
FDRSE #(.INIT(1'h0)) inst1 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[1]), .Q(inst1_Q));
FDRSE #(.INIT(1'h0)) inst2 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[2]), .Q(inst2_Q));
FDRSE #(.INIT(1'h0)) inst3 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[3]), .Q(inst3_Q));
FDRSE #(.INIT(1'h0)) inst4 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[4]), .Q(inst4_Q));
FDRSE #(.INIT(1'h0)) inst5 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[5]), .Q(inst5_Q));
FDRSE #(.INIT(1'h0)) inst6 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[6]), .Q(inst6_Q));
FDRSE #(.INIT(1'h0)) inst7 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[7]), .Q(inst7_Q));
FDRSE #(.INIT(1'h0)) inst8 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[8]), .Q(inst8_Q));
FDRSE #(.INIT(1'h0)) inst9 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[9]), .Q(inst9_Q));
FDRSE #(.INIT(1'h0)) inst10 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[10]), .Q(inst10_Q));
FDRSE #(.INIT(1'h0)) inst11 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[11]), .Q(inst11_Q));
FDRSE #(.INIT(1'h0)) inst12 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[12]), .Q(inst12_Q));
FDRSE #(.INIT(1'h0)) inst13 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[13]), .Q(inst13_Q));
FDRSE #(.INIT(1'h0)) inst14 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[14]), .Q(inst14_Q));
FDRSE #(.INIT(1'h0)) inst15 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[15]), .Q(inst15_Q));
FDRSE #(.INIT(1'h0)) inst16 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[16]), .Q(inst16_Q));
FDRSE #(.INIT(1'h0)) inst17 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[17]), .Q(inst17_Q));
FDRSE #(.INIT(1'h0)) inst18 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[18]), .Q(inst18_Q));
FDRSE #(.INIT(1'h0)) inst19 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[19]), .Q(inst19_Q));
FDRSE #(.INIT(1'h0)) inst20 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[20]), .Q(inst20_Q));
FDRSE #(.INIT(1'h0)) inst21 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[21]), .Q(inst21_Q));
FDRSE #(.INIT(1'h0)) inst22 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[22]), .Q(inst22_Q));
FDRSE #(.INIT(1'h0)) inst23 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[23]), .Q(inst23_Q));
FDRSE #(.INIT(1'h0)) inst24 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[24]), .Q(inst24_Q));
FDRSE #(.INIT(1'h0)) inst25 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[25]), .Q(inst25_Q));
FDRSE #(.INIT(1'h0)) inst26 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[26]), .Q(inst26_Q));
FDRSE #(.INIT(1'h0)) inst27 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[27]), .Q(inst27_Q));
FDRSE #(.INIT(1'h0)) inst28 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[28]), .Q(inst28_Q));
FDRSE #(.INIT(1'h0)) inst29 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[29]), .Q(inst29_Q));
FDRSE #(.INIT(1'h0)) inst30 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[30]), .Q(inst30_Q));
FDRSE #(.INIT(1'h0)) inst31 (.C(CLK), .CE(1'b1), .R(1'b0), .S(1'b0), .D(I[31]), .Q(inst31_Q));
assign O = {inst31_Q,inst30_Q,inst29_Q,inst28_Q,inst27_Q,inst26_Q,inst25_Q,inst24_Q,inst23_Q,inst22_Q,inst21_Q,inst20_Q,inst19_Q,inst18_Q,inst17_Q,inst16_Q,inst15_Q,inst14_Q,inst13_Q,inst12_Q,inst11_Q,inst10_Q,inst9_Q,inst8_Q,inst7_Q,inst6_Q,inst5_Q,inst4_Q,inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter32 (output [31:0] O, output  COUT, input  CLK);
wire [31:0] inst0_O;
wire  inst0_COUT;
wire [31:0] inst1_O;
Add32_cout inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register32 inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module main (output [7:0] LED, input  CLKIN);
wire [31:0] inst0_O;
wire  inst0_COUT;
Counter32 inst0 (.O(inst0_O), .COUT(inst0_COUT), .CLK(CLKIN));
assign LED = {inst0_O[31],inst0_O[30],inst0_O[29],inst0_O[28],inst0_O[27],inst0_O[26],inst0_O[25],inst0_O[24]};
endmodule

