module main (input [7:0] SWITCH, output [7:0] LED);
assign LED = SWITCH;
endmodule

