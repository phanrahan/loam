module FullAdder (input  I0, input  I1, input  CIN, output  O, output  COUT);
wire  inst0_O;
wire  inst1_CO;
SB_LUT4 #(.LUT_INIT(16'h9696)) inst0 (.I0(I0), .I1(I1), .I2(CIN), .I3(1'b0), .O(inst0_O));
SB_CARRY inst1 (.I0(I0), .I1(I1), .CI(CIN), .CO(inst1_CO));
assign O = inst0_O;
assign COUT = inst1_CO;
endmodule

module Add16Cout (input [15:0] I0, input [15:0] I1, output [15:0] O, output  COUT);
wire  inst0_O;
wire  inst0_COUT;
wire  inst1_O;
wire  inst1_COUT;
wire  inst2_O;
wire  inst2_COUT;
wire  inst3_O;
wire  inst3_COUT;
wire  inst4_O;
wire  inst4_COUT;
wire  inst5_O;
wire  inst5_COUT;
wire  inst6_O;
wire  inst6_COUT;
wire  inst7_O;
wire  inst7_COUT;
wire  inst8_O;
wire  inst8_COUT;
wire  inst9_O;
wire  inst9_COUT;
wire  inst10_O;
wire  inst10_COUT;
wire  inst11_O;
wire  inst11_COUT;
wire  inst12_O;
wire  inst12_COUT;
wire  inst13_O;
wire  inst13_COUT;
wire  inst14_O;
wire  inst14_COUT;
wire  inst15_O;
wire  inst15_COUT;
FullAdder inst0 (.I0(I0[0]), .I1(I1[0]), .CIN(1'b0), .O(inst0_O), .COUT(inst0_COUT));
FullAdder inst1 (.I0(I0[1]), .I1(I1[1]), .CIN(inst0_COUT), .O(inst1_O), .COUT(inst1_COUT));
FullAdder inst2 (.I0(I0[2]), .I1(I1[2]), .CIN(inst1_COUT), .O(inst2_O), .COUT(inst2_COUT));
FullAdder inst3 (.I0(I0[3]), .I1(I1[3]), .CIN(inst2_COUT), .O(inst3_O), .COUT(inst3_COUT));
FullAdder inst4 (.I0(I0[4]), .I1(I1[4]), .CIN(inst3_COUT), .O(inst4_O), .COUT(inst4_COUT));
FullAdder inst5 (.I0(I0[5]), .I1(I1[5]), .CIN(inst4_COUT), .O(inst5_O), .COUT(inst5_COUT));
FullAdder inst6 (.I0(I0[6]), .I1(I1[6]), .CIN(inst5_COUT), .O(inst6_O), .COUT(inst6_COUT));
FullAdder inst7 (.I0(I0[7]), .I1(I1[7]), .CIN(inst6_COUT), .O(inst7_O), .COUT(inst7_COUT));
FullAdder inst8 (.I0(I0[8]), .I1(I1[8]), .CIN(inst7_COUT), .O(inst8_O), .COUT(inst8_COUT));
FullAdder inst9 (.I0(I0[9]), .I1(I1[9]), .CIN(inst8_COUT), .O(inst9_O), .COUT(inst9_COUT));
FullAdder inst10 (.I0(I0[10]), .I1(I1[10]), .CIN(inst9_COUT), .O(inst10_O), .COUT(inst10_COUT));
FullAdder inst11 (.I0(I0[11]), .I1(I1[11]), .CIN(inst10_COUT), .O(inst11_O), .COUT(inst11_COUT));
FullAdder inst12 (.I0(I0[12]), .I1(I1[12]), .CIN(inst11_COUT), .O(inst12_O), .COUT(inst12_COUT));
FullAdder inst13 (.I0(I0[13]), .I1(I1[13]), .CIN(inst12_COUT), .O(inst13_O), .COUT(inst13_COUT));
FullAdder inst14 (.I0(I0[14]), .I1(I1[14]), .CIN(inst13_COUT), .O(inst14_O), .COUT(inst14_COUT));
FullAdder inst15 (.I0(I0[15]), .I1(I1[15]), .CIN(inst14_COUT), .O(inst15_O), .COUT(inst15_COUT));
assign O = {inst15_O,inst14_O,inst13_O,inst12_O,inst11_O,inst10_O,inst9_O,inst8_O,inst7_O,inst6_O,inst5_O,inst4_O,inst3_O,inst2_O,inst1_O,inst0_O};
assign COUT = inst15_COUT;
endmodule

module Register16 (input [15:0] I, output [15:0] O, input  CLK);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
wire  inst4_Q;
wire  inst5_Q;
wire  inst6_Q;
wire  inst7_Q;
wire  inst8_Q;
wire  inst9_Q;
wire  inst10_Q;
wire  inst11_Q;
wire  inst12_Q;
wire  inst13_Q;
wire  inst14_Q;
wire  inst15_Q;
SB_DFF inst0 (.C(CLK), .D(I[0]), .Q(inst0_Q));
SB_DFF inst1 (.C(CLK), .D(I[1]), .Q(inst1_Q));
SB_DFF inst2 (.C(CLK), .D(I[2]), .Q(inst2_Q));
SB_DFF inst3 (.C(CLK), .D(I[3]), .Q(inst3_Q));
SB_DFF inst4 (.C(CLK), .D(I[4]), .Q(inst4_Q));
SB_DFF inst5 (.C(CLK), .D(I[5]), .Q(inst5_Q));
SB_DFF inst6 (.C(CLK), .D(I[6]), .Q(inst6_Q));
SB_DFF inst7 (.C(CLK), .D(I[7]), .Q(inst7_Q));
SB_DFF inst8 (.C(CLK), .D(I[8]), .Q(inst8_Q));
SB_DFF inst9 (.C(CLK), .D(I[9]), .Q(inst9_Q));
SB_DFF inst10 (.C(CLK), .D(I[10]), .Q(inst10_Q));
SB_DFF inst11 (.C(CLK), .D(I[11]), .Q(inst11_Q));
SB_DFF inst12 (.C(CLK), .D(I[12]), .Q(inst12_Q));
SB_DFF inst13 (.C(CLK), .D(I[13]), .Q(inst13_Q));
SB_DFF inst14 (.C(CLK), .D(I[14]), .Q(inst14_Q));
SB_DFF inst15 (.C(CLK), .D(I[15]), .Q(inst15_Q));
assign O = {inst15_Q,inst14_Q,inst13_Q,inst12_Q,inst11_Q,inst10_Q,inst9_Q,inst8_Q,inst7_Q,inst6_Q,inst5_Q,inst4_Q,inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter16 (output [15:0] O, output  COUT, input  CLK);
wire [15:0] inst0_O;
wire  inst0_COUT;
wire [15:0] inst1_O;
Add16Cout inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register16 inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module And2 (input [1:0] I, output  O);
wire  inst0_O;
SB_LUT4 #(.LUT_INIT(16'h8888)) inst0 (.I0(I[0]), .I1(I[1]), .I2(1'b0), .I3(1'b0), .O(inst0_O));
assign O = inst0_O;
endmodule

module Mux2 (input [1:0] I, input  S, output  O);
wire  inst0_O;
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst0 (.I0(I[0]), .I1(I[1]), .I2(S), .I3(1'b0), .O(inst0_O));
assign O = inst0_O;
endmodule

module main (input [4:0] J1, output [3:0] J3, input  CLKIN);
wire [15:0] inst0_O;
wire  inst0_COUT;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_O;
wire  inst4_Q;
wire  inst5_O;
wire  inst6_Q;
wire  inst7_O;
wire  inst8_O;
wire  inst9_Q;
wire  inst10_Q;
wire  inst11_Q;
wire  inst12_O;
wire  inst13_O;
wire  inst14_O;
wire  inst15_O;
wire  inst16_O;
wire  inst17_O;
wire  inst18_O;
wire  inst19_O;
wire  inst20_O;
wire  inst21_O;
wire  inst22_O;
wire  inst23_O;
Counter16 inst0 (.O(inst0_O), .COUT(inst0_COUT), .CLK(CLKIN));
SB_DFFE inst1 (.C(CLKIN), .E(inst0_COUT), .D(J1[4]), .Q(inst1_Q));
SB_DFFE inst2 (.C(CLKIN), .E(inst0_COUT), .D(inst1_Q), .Q(inst2_Q));
And2 inst3 (.I({inst2_Q,inst1_Q}), .O(inst3_O));
SB_DFF inst4 (.C(CLKIN), .D(inst3_O), .Q(inst4_Q));
SB_LUT4 #(.LUT_INIT(16'h4444)) inst5 (.I0(inst3_O), .I1(inst4_Q), .I2(1'b0), .I3(1'b0), .O(inst5_O));
SB_DFFE inst6 (.C(CLKIN), .E(inst5_O), .D(inst7_O), .Q(inst6_Q));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst7 (.I0(inst14_O), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst7_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst8 (.I0(inst6_Q), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst8_O));
SB_DFFE inst9 (.C(CLKIN), .E(inst5_O), .D(inst17_O), .Q(inst9_Q));
SB_DFFE inst10 (.C(CLKIN), .E(inst5_O), .D(inst20_O), .Q(inst10_Q));
SB_DFFE inst11 (.C(CLKIN), .E(inst5_O), .D(inst23_O), .Q(inst11_Q));
SB_LUT4 #(.LUT_INIT(16'hF888)) inst12 (.I0(inst10_Q), .I1(J1[0]), .I2(inst11_Q), .I3(J1[0]), .O(inst12_O));
SB_LUT4 #(.LUT_INIT(16'h0001)) inst13 (.I0(J1[1]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst13_O));
Mux2 inst14 (.I({inst13_O,inst12_O}), .S(inst8_O), .O(inst14_O));
SB_LUT4 #(.LUT_INIT(16'hF888)) inst15 (.I0(inst8_O), .I1(J1[1]), .I2(1'b0), .I3(1'b0), .O(inst15_O));
SB_LUT4 #(.LUT_INIT(16'h0001)) inst16 (.I0(J1[2]), .I1(J1[3]), .I2(1'b0), .I3(1'b0), .O(inst16_O));
Mux2 inst17 (.I({inst16_O,inst15_O}), .S(inst9_Q), .O(inst17_O));
SB_LUT4 #(.LUT_INIT(16'hF888)) inst18 (.I0(inst9_Q), .I1(J1[2]), .I2(1'b0), .I3(1'b0), .O(inst18_O));
SB_LUT4 #(.LUT_INIT(16'h0001)) inst19 (.I0(J1[3]), .I1(J1[0]), .I2(1'b0), .I3(1'b0), .O(inst19_O));
Mux2 inst20 (.I({inst19_O,inst18_O}), .S(inst10_Q), .O(inst20_O));
SB_LUT4 #(.LUT_INIT(16'hF888)) inst21 (.I0(inst9_Q), .I1(J1[3]), .I2(inst10_Q), .I3(J1[3]), .O(inst21_O));
SB_LUT4 #(.LUT_INIT(16'h0001)) inst22 (.I0(J1[0]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst22_O));
Mux2 inst23 (.I({inst22_O,inst21_O}), .S(inst11_Q), .O(inst23_O));
assign J3 = {inst11_Q,inst10_Q,inst9_Q,inst8_O};
endmodule

