module main (output  D1, output  D2, output  D3, output  D4);
assign D1 = 1'b1;
assign D2 = 1'b1;
assign D3 = 1'b1;
assign D4 = 1'b1;
endmodule

