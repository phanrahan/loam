module main (output  LED1, output  LED2);
assign LED1 = 1'b1;
assign LED2 = 1'b1;
endmodule

