module main (input  S2, input  S4, input  S1, input  S3, output  D1, output  D2, output  D3, output  D4);
assign D1 = S1;
assign D2 = S2;
assign D3 = S3;
assign D4 = S4;
endmodule

