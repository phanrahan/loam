module main (output  LED1, input  RST_N);
assign LED1 = RST_N;
endmodule

