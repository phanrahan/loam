module main (output  PIN2);
assign PIN2 = 1'b1;
endmodule

