module main (output  LED);
assign LED = 1'b1;
endmodule

